module ID_EX_reg (nextPC ,ReadData1 ,ReadData2 ,signExtendResult ,);




endmodule
