module ForwardingUnit();




endmodule
